library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity Mux_we is
    port (
      D : in std_logic_vector(0 to 3);
      sel : in std_logic_vector(0 to 1);
      y : out std_logic
    ) ;
  end Mux_we ;

architecture Mux_arch_when_else of Mux_we is
begin
  y <=  D(0) when sel = "00" else
        D(1) when sel = "01" else
        D(2) when sel = "10" else
        D(3) when sel = "11" else
        '0';
end Mux_arch_when_else ;